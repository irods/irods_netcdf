  netcdf example {   // example of CDL notation
  dimensions:
          time = 20;
          depth = 3;
	  lon = 3 ;
	  lat = 40 ;
  variables:
	  float rh(lon, lat) ; // lon, lat
		  rh:units = "percent" ;
		  rh:long_name = "Relative humidity" ;
  // global attributes
	  :title = "Simple example, lacks some conventions" ;
  data:


   rh =
  2.1, 3.1, 5.1, 7.1, 11.1, 13.1, 17.1, 19.1,
  2.3, 3.3, 5.3, 7.3, 11.3, 13.3, 17.3, 19.3,
  2.5, 3.5, 5.5, 7.5, 11.5, 13.5, 17.5, 19.5,
  2.7, 3.7, 5.7, 7.7, 11.7, 13.7, 17.7, 19.7,
  2.9, 3.9, 5.9, 7.9, 11.9, 13.9, 17.9, 19.9,

  23.1, 29.1, 31.1, 37.1, 41.1, 43.1, 47.1, 53.1,
  23.3, 29.3, 31.3, 37.3, 41.3, 43.3, 47.3, 53.3,
  23.5, 29.5, 31.5, 37.5, 41.5, 43.5, 47.5, 53.5,
  23.7, 29.7, 31.7, 37.7, 41.7, 43.7, 47.7, 53.7,
  23.9, 29.9, 31.9, 37.9, 41.9, 43.9, 47.9, 53.9,

   59.1, 61.1, 67.1, 71.1, 73.1, 79.1, 83.1, 89.1,
   59.3, 61.3, 67.3, 71.3, 73.3, 79.3, 83.3, 89.3,
   59.5, 61.5, 67.5, 71.5, 73.5, 79.5, 83.5, 89.5,
   59.7, 61.7, 67.7, 71.7, 73.7, 79.7, 83.7, 89.7,
   59.9, 61.9, 67.9, 71.9, 73.9, 79.9, 83.9, 89.9;

  }
//time[10:1:12] depth[3:1:3] lat[4:1:7] lon[30:1:34]
